/**
 * 1-bit register:
 * If load[t] == 1 then out[t+1] = in[t]
 *    else out does not change (out[t+1] = out[t])
 */

`default_nettype none
module Bit(
	input clk,
	input in,
	input load,
	output out
);


	//..LET THE DRAMA begin
	// //USING MUX AND DFF
	// Mux PICK(
	// 	// in,
	// );

	reg bit_out;
	reg	load_out;
	always @(posedge clk) begin
		if (load)
		bit_out <= in;
	end

	assign out = bit_out;
endmodule
